entity audio_and_video_config is (
	port(
		clock_50;
		reset,
		
		i2c_sdat,
		i2c_sclk
	);
)

generic 